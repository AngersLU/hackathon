`define INDEX_32  1'b1
`define INDEX    32